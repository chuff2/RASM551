`timescale 100ps / 10ps
module LA_dig_tb();
 parameter ENTRIES = 384,	// defaults to 384 for simulation, use 12288 for DE-0
            LOG2 = 9;		// Log base 2 of number of entries
			
			
localparam TRIG_CFG_WR = {2'b01, 6'h0};
localparam TRIG_CFG_RD = {2'b00, 6'h0};
	
localparam CH1TrigCfgWr = {2'b01, 6'h01};
localparam CH2TrigCfgWr = {2'b01, 6'h02};
localparam CH3TrigCfgWr = {2'b01, 6'h03};
localparam CH4TrigCfgWr = {2'b01, 6'h04};
localparam CH5TrigCfgWr = {2'b01, 6'h05};
	
localparam CH1TrigCfgRd = {2'b0, 6'h01};
localparam CH2TrigCfgRd = {2'b0, 6'h02};
localparam CH3TrigCfgRd = {2'b0, 6'h03};
localparam CH4TrigCfgRd = {2'b0, 6'h04};
localparam CH5TrigCfgRd = {2'b0, 6'h05};
	
//// Interconnects to DUT/support defined as type wire /////
wire clk400MHz,locked;			// PLL output signals to DUT
wire clk;						// 100MHz clock generated at this level from clk400MHz
wire VIH_PWM,VIL_PWM;			// connect to PWM outputs to monitor
logic CH1L,CH1H,CH2L,CH2H,CH3L;	// channel data inputs from AFE model
logic CH3H,CH4L,CH4H,CH5L,CH5H;	// channel data inputs from AFE model
wire RX,TX;						// interface to host
wire cmd_sent,resp_rdy;			// from master UART, monitored in test bench
wire [7:0] resp;				// from master UART, reponse received from DUT
wire tx_prot;					// UART signal for protocol triggering
wire SS_n,SCLK,MOSI;			// SPI signals for SPI protocol triggering
wire CH1L_mux,CH1H_mux;         // output of muxing logic for CH1 to enable testing of protocol triggering
wire CH2L_mux,CH2H_mux;			// output of muxing logic for CH2 to enable testing of protocol triggering
wire CH3L_mux,CH3H_mux;			// output of muxing logic for CH3 to enable testing of protocol triggering

////// Stimulus is declared as type reg ///////
reg REF_CLK, RST_n;
reg [15:0] host_cmd;			// command host is sending to DUT
reg send_cmd;					// asserted to initiate sending of command
reg clr_resp_rdy;				// asserted to knock down resp_rdy
reg [1:0] clk_div;				// counter used to derive 100MHz clk from clk400MHz
reg strt_tx;					// kick off unit used for protocol triggering

logic UART_triggering;
logic SPI_triggering;

/////////////////////////////////////////////////////////////
// Channel Dumps can be written to file to aid in testing //
///////////////////////////////////////////////////////////
// setup file pointers here if going to do that

///////////////////////////
// Define command bytes //
/////////////////////////
// May or may not want to make some localparams to represent command bytes to LA core
localparam READ = 2'b00;
localparam WRITE = 2'b01;
localparam DUMP = 2'b10;

/////////////////////////////////
// localparam UART_triggering = 1'b0;	// set to true if testing UART based triggering
// localparam SPI_triggering = 1'b1;	// set to true if testing SPI based triggering
// UART and SPI triggering is based off the TrigCfg register
assign UART_triggering = ~iDUT.iDIG.TrigCfg[0];
assign SPI_triggering = ~iDUT.iDIG.TrigCfg[1];


///// Instantiate Analog Front End model (provides stimulus to channels) ///////
AFE iAFE(.smpl_clk(clk400MHz),.VIH_PWM(VIH_PWM),.VIL_PWM(VIL_PWM),
         .CH1L(CH1L),.CH1H(CH1H),.CH2L(CH2L),.CH2H(CH2H),.CH3L(CH3L),
         .CH3H(CH3H),.CH4L(CH4L),.CH4H(CH4H),.CH5L(CH5L),.CH5H(CH5H));
		 
//// Mux for muxing in protocol triggering for CH1 /////
assign {CH1H_mux,CH1L_mux} = (UART_triggering) ? {2{tx_prot}} :		// assign to output of UART_tx used to test UART triggering
                             (SPI_triggering) ? {2{SS_n}}: 			// assign to output of SPI SS_n if SPI triggering
				             {CH1H,CH1L};

//// Mux for muxing in protocol triggering for CH2 /////
assign {CH2H_mux,CH2L_mux} = (SPI_triggering) ? {2{SCLK}}: 			// assign to output of SPI SCLK if SPI triggering
				             {CH2H,CH2L};	

//// Mux for muxing in protocol triggering for CH3 /////
assign {CH3H_mux,CH3L_mux} = (SPI_triggering) ? {2{MOSI}}: 			// assign to output of SPI MOSI if SPI triggering
				             {CH3H,CH3L};					  
	 
////// Instantiate DUT //////// TODO do we need the LED?? It wasnt in there originally but I added it in to get rid of error
LA_dig iDUT(.clk400MHz(clk400MHz),.RST_n(RST_n),.locked(locked),
            .VIH_PWM(VIH_PWM),.VIL_PWM(VIL_PWM),.CH1L(CH1L_mux),.CH1H(CH1H_mux),
			.CH2L(CH2L_mux),.CH2H(CH2H_mux),.CH3L(CH3L_mux),.CH3H(CH3H_mux),.CH4L(CH4L),
			.CH4H(CH4H),.CH5L(CH5L),.CH5H(CH5H),.RX(RX),.TX(TX), .LED());



///// Instantiate PLL to provide 400MHz clk from 50MHz ///////
pll8x iPLL(.ref_clk(REF_CLK),.RST_n(RST_n),.out_clk(clk400MHz),.locked(locked));

///// It is useful to have a 100MHz clock at this level similar //////
///// to main system clock (clk).  So we will create one        //////
always @(posedge clk400MHz, negedge locked)
  if (~locked)
    clk_div <= 2'b00;
  else
    clk_div <= clk_div+1;
assign clk = clk_div[1];

//// Instantiate Master UART (mimics host commands) //////
/* unmodified version 
UART_comm_mstr iMSTR(.clk(clk), .rst_n(RST_n), .RX(TX), .TX(RX),
                     .cmd(host_cmd), .send_cmd(send_cmd),
					 .cmd_sent(cmd_sent), .resp_rdy(resp_rdy),
					 .resp(resp), .clr_resp_rdy(clr_resp_rdy));
*/
CommMaster iMSTR(.clk(clk), .rst_n(RST_n), .RX(TX), .TX(RX),
                     .cmd(host_cmd), .snd_cmd(send_cmd),
					 .cmd_cmplt(cmd_sent), .resp_cmplt(resp_rdy),
					 .resp(resp), .clr_rdy(clr_resp_rdy));
					 
////////////////////////////////////////////////////////////////
// Instantiate transmitter as source for protocol triggering //
//////////////////////////////////////////////////////////////
/* unmodified version
uart_tx iTX(.clk(clk), .rst_n(RST_n), .tx(tx_prot), .strt_tx(strt_tx),
        .tx_data(8'h96), .tx_done());
*/
uart_tx iTX(.clk(clk), .rst_n(RST_n), .TX(tx_prot), .trmt(strt_tx),
        .tx_data(8'h96), .tx_done());

					 
////////////////////////////////////////////////////////////////////
// Instantiate SPI transmitter as source for protocol triggering //
//////////////////////////////////////////////////////////////////
SPI_mstr iSPI(.clk(clk),.rst_n(RST_n),.SS_n(SS_n),.SCLK(SCLK),.wrt(strt_tx),.done(done),
              .data_out(16'h6600),.MOSI(MOSI),.pos_edge(1'b0),.width8(1'b1));


/********************************************************************
* Signals for chan_trig_test
********************************************************************/
logic [10:0] channels;
logic [5:0] CHTrigCfg;
logic [9:0] prevChannels;
		
logic [7:0] dataRead;
logic error;

initial begin
//   put your testing code here.
REF_CLK = 0;
RST_n = 0;
host_cmd = 16'h0000;//read address 0			
send_cmd = 0;					
clr_resp_rdy = 0;				
clk_div = 0;				
strt_tx = 0;	

repeat(3) @(negedge clk)
RST_n = 1;
strt_tx = 1;
send_cmd = 1;
@(negedge clk) send_cmd = 0;

repeat (10) @(negedge clk);
// test1();
//test2();
//test4(4'h1, 8'h86);
//test5;
chan_trig_test;
$stop;
end

always
  #100 REF_CLK = ~REF_CLK;

///// Perhaps put some basic tasks in a separate file to keep your test bench less cluttered /////
`include "tb_tasks.sv"
`include "test1.sv";
`include "test2.sv";
`include "test4.sv";
`include "test5.sv";
`include "chan_trig_test.sv";

endmodule	
