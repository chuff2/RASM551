module prot_trig();





endmodule
